
module IF_Stage(clk, rst, 