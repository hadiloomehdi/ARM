`timescale 1ns/1ns
module Controller(output reg Flush,Branch_Taken );
  
  assign {Flush,Branch_Taken} =  2'b0;

endmodule
